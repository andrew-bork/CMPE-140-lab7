module regfile (
        input  wire        clk,
        input  wire        we,
        input  wire [4:0]  ra1,
        input  wire [4:0]  ra2,
        input  wire [4:0]  ra3,
        input  wire [4:0]  wa,
        input  wire [31:0] wd,
        output wire [31:0] rd1,
        output wire [31:0] rd2,
        output wire [31:0] rd3
    );

    reg [31:0] rf [0:31];

    integer n;
    
    initial begin
        for (n = 0; n < 32; n = n + 1) rf[n] = 32'h0;
        rf[29] = 32'h100; // Initialze $sp
    end
    
    always @ (posedge clk) begin
        if (we) rf[wa] <= wd;
    end

    assign rd1 = (ra1 == 0) ? 0 : rf[ra1];
    assign rd2 = (ra2 == 0) ? 0 : rf[ra2];
    assign rd3 = (ra3 == 0) ? 0 : rf[ra3];

    
    initial begin
        $dumpfile("mips.vcd");
        $dumpvars(0, rf[7]);
        $dumpvars(0, rf[8]);
        $dumpvars(0, rf[3]);
        $dumpvars(0, rf[31]);
        $dumpvars(0, rf[16]);
        $dumpvars(0, rf[4]);
        $dumpvars(0, rf[2]);
        $dumpvars(0, rf[29]);
    end

endmodule